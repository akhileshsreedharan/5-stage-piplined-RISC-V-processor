//opcodes
`define RV32_BRANCH 7'b1100011
`define RV32_JAL    7'b1101111
`define RV32_LOAD   7'b0000011
`define RV32_STORE  7'b0100011
`define RV32_RTYPE  7'b0110011
`define RV32_OP_IMM 7'b0010011

//funct3 encoding
`define RV32_FUNCT3_BRANCH_BEQ  3'b000
`define RV32_FUNCT3_BRANCH_BNE  3'b001
`define RV32_FUNCT3_BRANCH_BLT  3'b100
`define RV32_FUNCT3_BRANCH_BGE  3'b101
`define RV32_FUNCT3_BRANCH_BLTU 3'b110
`define RV32_FUNCT3_BRANCH_BGEU 3'b111



`define RV32_FUNCT3_LOAD       3'b011

`define RV32_FUNCT3_STORE      3'b111

`define RV32_FUNCT3_ADDI       3'b000
`define RV32_FUNCT3_SLLI       3'b001
`define RV32_FUNCT3_SRLI       3'b101

`define RV32_FUNCT3_RTYPE_ADD  3'b000
`define RV32_FUNCT3_RTYPE_SUB  3'b000
`define RV32_FUNCT3_RTYPE_SLL  3'b001
`define RV32_FUNCT3_RTYPE_XOR  3'b100
//`define RV32_FUNCT3_RTYPE_SRL  3'b101
//`define RV32_FUNCT3_RTYPE_SRA  3'b101
`define RV32_FUNCT3_RTYPE_OR   3'b110
`define RV32_FUNCT3_RTYPE_AND  3'b111

`define RV32_FUNCT3_RTYPE_INVALID  3'b010


//funct7 encoding
`define RV32_FUNCT7_RTYPE_ADD  7'b0000000
`define RV32_FUNCT7_RTYPE_SUB  7'b0100000
//`define RV32_FUNCT7_RTYPE_SLL  7'b0000000
`define RV32_FUNCT7_RTYPE_XOR  7'b0000000
//`define RV32_FUNCT7_RTYPE_SRL  7'b0000000
//`define RV32_FUNCT7_RTYPE_SRA  7'b0100000
`define RV32_FUNCT7_RTYPE_OR   7'b0000000
`define RV32_FUNCT7_RTYPE_AND  7'b0000000
`define RV32_FUNCT7_RTYPE_INVALID  7'b1111111

`define RV32_FUNCT7_RTYPE_SLLI  7'b0000000
`define RV32_FUNCT7_RTYPE_SRLI  7'b0000000
